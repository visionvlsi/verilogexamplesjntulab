module fa(a,b,cin,sum,co);
input a,b,cin;
output sum,co;
ha ha1(a,b,s1,c1);
ha ha2(cin,s1,sum,c2);
or or1(co,c1,c2);
endmodule
